`timescale 1ns / 1ps

module systolic_matrix_mult_3x3_tb;
    
    // Parameters for 3x3 matrices
    parameter DATA_WIDTH = 16;
    parameter FRAC_WIDTH = 8;
    parameter M = 3;  // Rows of A, rows of C
    parameter N = 3;  // Cols of B, cols of C
    parameter K = 3;  // Cols of A, rows of B
    
    // DUT signals
    reg clk;
    reg rst_n;
    reg start;
    
    // Matrix A input
    reg signed [DATA_WIDTH-1:0] a_data;
    reg [$clog2(M)-1:0] a_row;
    reg [$clog2(K)-1:0] a_col;
    reg a_valid;
    
    // Matrix B input
    reg signed [DATA_WIDTH-1:0] b_data;
    reg [$clog2(K)-1:0] b_row;
    reg [$clog2(N)-1:0] b_col;
    reg b_valid;
    
    // Matrix C output
    wire signed [DATA_WIDTH-1:0] c_data;
    wire [$clog2(M)-1:0] c_row;
    wire [$clog2(N)-1:0] c_col;
    wire c_valid;
    wire done;
    
    // Test storage
    reg signed [DATA_WIDTH-1:0] test_a [0:M-1][0:K-1];
    reg signed [DATA_WIDTH-1:0] test_b [0:K-1][0:N-1];
    reg signed [DATA_WIDTH-1:0] expected_c [0:M-1][0:N-1];
    reg signed [DATA_WIDTH-1:0] result_c [0:M-1][0:N-1];
    
    // Instantiate DUT - using v2 which has better control logic
    systolic_matrix_mult #(
        .DATA_WIDTH(DATA_WIDTH),
        .FRAC_WIDTH(FRAC_WIDTH),
        .M(M),
        .N(N),
        .K(K)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .start(start),
        .a_data(a_data),
        .a_row(a_row),
        .a_col(a_col),
        .a_valid(a_valid),
        .b_data(b_data),
        .b_row(b_row),
        .b_col(b_col),
        .b_valid(b_valid),
        .c_data(c_data),
        .c_row(c_row),
        .c_col(c_col),
        .c_valid(c_valid),
        .done(done)
    );
    
    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    // Fixed-point conversion functions
    function signed [DATA_WIDTH-1:0] to_fixed(input real val);
        begin
            to_fixed = val * (1 << FRAC_WIDTH);
        end
    endfunction
    
    function real from_fixed(input signed [DATA_WIDTH-1:0] val);
        begin
            from_fixed = $itor(val) / (1 << FRAC_WIDTH);
        end
    endfunction
    
    // Test tasks
    integer i, j, k;
    
    // Initialize test case
    task init_test_case;
        begin
            $display("\nTest: 3x3 Systolic Array Matrix Multiplication");
            $display("\nTest Case 1: Simple Sequential Pattern");
            // Matrix A: Sequential values 1-9
            test_a[0][0] = to_fixed(1.0); test_a[0][1] = to_fixed(2.0); test_a[0][2] = to_fixed(3.0);
            test_a[1][0] = to_fixed(4.0); test_a[1][1] = to_fixed(5.0); test_a[1][2] = to_fixed(6.0);
            test_a[2][0] = to_fixed(7.0); test_a[2][1] = to_fixed(8.0); test_a[2][2] = to_fixed(9.0);
            
            // Matrix B: Identity matrix (should return A)
            test_b[0][0] = to_fixed(1.0); test_b[0][1] = to_fixed(0.0); test_b[0][2] = to_fixed(0.0);
            test_b[1][0] = to_fixed(0.0); test_b[1][1] = to_fixed(1.0); test_b[1][2] = to_fixed(0.0);
            test_b[2][0] = to_fixed(0.0); test_b[2][1] = to_fixed(0.0); test_b[2][2] = to_fixed(1.0);
            
            $display("Matrix A:");
            for (i = 0; i < M; i = i + 1) begin
                $write("  [");
                for (j = 0; j < K; j = j + 1) begin
                    $write("%6.1f ", from_fixed(test_a[i][j]));
                end
                $display("]");
            end
            
            $display("Matrix B (Identity):");
            for (i = 0; i < K; i = i + 1) begin
                $write("  [");
                for (j = 0; j < N; j = j + 1) begin
                    $write("%6.1f ", from_fixed(test_b[i][j]));
                end
                $display("]");
            end
        end
    endtask
    
    // Initialize second test case
    task init_test_case_2;
        begin
            $display("\nTest Case 2: Non-trivial Multiplication");
            // Matrix A
            test_a[0][0] = to_fixed(2.0); test_a[0][1] = to_fixed(1.0); test_a[0][2] = to_fixed(3.0);
            test_a[1][0] = to_fixed(1.0); test_a[1][1] = to_fixed(4.0); test_a[1][2] = to_fixed(2.0);
            test_a[2][0] = to_fixed(3.0); test_a[2][1] = to_fixed(2.0); test_a[2][2] = to_fixed(1.0);
            
            // Matrix B
            test_b[0][0] = to_fixed(1.0); test_b[0][1] = to_fixed(2.0); test_b[0][2] = to_fixed(1.0);
            test_b[1][0] = to_fixed(3.0); test_b[1][1] = to_fixed(1.0); test_b[1][2] = to_fixed(2.0);
            test_b[2][0] = to_fixed(2.0); test_b[2][1] = to_fixed(1.0); test_b[2][2] = to_fixed(3.0);
            
            $display("Matrix A:");
            for (i = 0; i < M; i = i + 1) begin
                $write("  [");
                for (j = 0; j < K; j = j + 1) begin
                    $write("%6.1f ", from_fixed(test_a[i][j]));
                end
                $display("]");
            end
            
            $display("Matrix B:");
            for (i = 0; i < K; i = i + 1) begin
                $write("  [");
                for (j = 0; j < N; j = j + 1) begin
                    $write("%6.1f ", from_fixed(test_b[i][j]));
                end
                $display("]");
            end
        end
    endtask
    
    // Compute expected result
    task compute_expected;
        reg signed [2*DATA_WIDTH-1:0] temp_sum;
        begin
            for (i = 0; i < M; i = i + 1) begin
                for (j = 0; j < N; j = j + 1) begin
                    temp_sum = 0;
                    for (k = 0; k < K; k = k + 1) begin
                        temp_sum = temp_sum + (test_a[i][k] * test_b[k][j]);
                    end
                    expected_c[i][j] = temp_sum[DATA_WIDTH+FRAC_WIDTH-1:FRAC_WIDTH];
                end
            end
            
            // Display expected results
            $display("Expected Matrix C:");
            for (i = 0; i < M; i = i + 1) begin
                $write("  [");
                for (j = 0; j < N; j = j + 1) begin
                    $write("%6.1f ", from_fixed(expected_c[i][j]));
                end
                $display("]");
            end
        end
    endtask
    
    // Load matrix A into DUT
    task load_matrix_a;
        integer a_i, a_j;
        begin
            for (a_i = 0; a_i < M; a_i = a_i + 1) begin
                for (a_j = 0; a_j < K; a_j = a_j + 1) begin
                    @(posedge clk);
                    a_data = test_a[a_i][a_j];
                    a_row = a_i;
                    a_col = a_j;
                    a_valid = 1;
                end
            end
            @(posedge clk);
            a_valid = 0;
        end
    endtask
    
    // Load matrix B into DUT
    task load_matrix_b;
        integer b_i, b_j;
        begin
            for (b_i = 0; b_i < K; b_i = b_i + 1) begin
                for (b_j = 0; b_j < N; b_j = b_j + 1) begin
                    @(posedge clk);
                    b_data = test_b[b_i][b_j];
                    b_row = b_i;
                    b_col = b_j;
                    b_valid = 1;
                end
            end
            @(posedge clk);
            b_valid = 0;
        end
    endtask
    
    // Collect output matrix C
    task collect_result;
        begin
            // Initialize result matrix
            for (i = 0; i < M; i = i + 1) begin
                for (j = 0; j < N; j = j + 1) begin
                    result_c[i][j] = 0;
                end
            end
            
            while (!done) begin
                @(posedge clk);
                if (c_valid) begin
                    result_c[c_row][c_col] = c_data;
                    $display("Output C[%0d][%0d] = %f", c_row, c_col, from_fixed(c_data));
                end
            end
        end
    endtask
    
    // Compare results
    task check_results;
        reg test_passed;
        begin
            test_passed = 1;
            $display("\nComparing results:");
            for (i = 0; i < M; i = i + 1) begin
                for (j = 0; j < N; j = j + 1) begin
                    if (result_c[i][j] == expected_c[i][j]) begin
                        $display("PASS: C[%0d][%0d] = %f", i, j, from_fixed(result_c[i][j]));
                    end else begin
                        $display("FAIL: C[%0d][%0d] = %f (expected %f)", 
                            i, j, from_fixed(result_c[i][j]), from_fixed(expected_c[i][j]));
                        test_passed = 0;
                    end
                end
            end
            
            if (test_passed)
                $display("Test PASSED!");
            else
                $display("Test FAILED!");
        end
    endtask
    
    // Run a complete test
    task run_test;
        begin
            compute_expected();
            
            // Reset
            @(posedge clk);
            rst_n = 0;
            @(posedge clk);
            @(posedge clk);
            rst_n = 1;
            @(posedge clk);
            
            // Start operation
            start = 1;
            @(posedge clk);
            start = 0;
            
            // Load matrices in parallel
            fork
                load_matrix_a();
                load_matrix_b();
            join
            
            // Wait for computation and collect results
            collect_result();
            
            // Check results
            check_results();
            
            // Display timing information
            $display("\nSystolic array (3x3) completed in %0d cycles", 
                (M + N + K - 1));
            $display("Expected: %0d cycles for systolic operation", M + N + K - 1);
            $display("Sequential would take: %0d cycles", M * N * K);
        end
    endtask
    
    // Main test
    initial begin
        // Generate VCD for debugging
        $dumpfile("systolic_matrix_mult_3x3_tb.vcd");
        $dumpvars(0, systolic_matrix_mult_3x3_tb);
        
        // Initialize
        rst_n = 0;
        start = 0;
        a_valid = 0;
        b_valid = 0;
        
        // Run Test Case 1: Identity multiplication
        $display("\n======== TEST CASE 1: Identity Matrix Multiplication ========");
        init_test_case();
        run_test();
        
        #100;
        
        // Run Test Case 2: General multiplication
        $display("\n\n======== TEST CASE 2: General Matrix Multiplication ========");
        init_test_case_2();
        run_test();
        
        #100;
        $display("\n======== All 3x3 Tests Completed ========");
        $finish;
    end
    
    // Timeout watchdog
    initial begin
        #100000;
        $display("ERROR: Test timeout!");
        $finish;
    end

endmodule